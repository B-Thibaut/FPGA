-- Copyright (C) 2023  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 23.1std.0 Build 991 11/28/2023 SC Lite Edition"
-- CREATED		"Mon Apr 22 10:37:23 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY full_adder_4b IS 
	PORT
	(
		Cin :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		A2 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		A3 :  IN  STD_LOGIC;
		B4 :  IN  STD_LOGIC;
		A4 :  IN  STD_LOGIC;
		S1 :  OUT  STD_LOGIC;
		S2 :  OUT  STD_LOGIC;
		S3 :  OUT  STD_LOGIC;
		S4 :  OUT  STD_LOGIC;
		C :  OUT  STD_LOGIC
	);
END full_adder_4b;

ARCHITECTURE bdf_type OF full_adder_4b IS 

COMPONENT full_adder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 cin : IN STD_LOGIC;
		 Sum : OUT STD_LOGIC;
		 Cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;


BEGIN 



b2v_inst : full_adder
PORT MAP(A => A1,
		 B => B1,
		 cin => Cin,
		 Sum => S1,
		 Cout => SYNTHESIZED_WIRE_0);


b2v_inst1 : full_adder
PORT MAP(A => A2,
		 B => B2,
		 cin => SYNTHESIZED_WIRE_0,
		 Sum => S2,
		 Cout => SYNTHESIZED_WIRE_1);


b2v_inst2 : full_adder
PORT MAP(A => A3,
		 B => B3,
		 cin => SYNTHESIZED_WIRE_1,
		 Sum => S3,
		 Cout => SYNTHESIZED_WIRE_2);


b2v_inst3 : full_adder
PORT MAP(A => A4,
		 B => B4,
		 cin => SYNTHESIZED_WIRE_2,
		 Sum => S4,
		 Cout => C);


END bdf_type;